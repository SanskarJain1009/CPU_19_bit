//Logic for Adder

module adder(
input [18:0] a,b,
output [18:0] sum
);
assign sum = a + b;
endmodule
